module MyNameROM(
	input VGA_CLK,
	input [5:0] address,
	output reg [63:0] data
);
always @(posedge VGA_CLK)
	begin
	case(address)
	//Ahmad
	00: data <= 64'd0000000000000000000;
	01: data <= 64'd0000000000000000000;
	02: data <= 64'd0000000072477573148;
	03: data <= 64'd0000000242128781324;
	04: data <= 64'd0000000465467080716;
	05: data <= 64'd0000000852230552636;
	06: data <= 64'd0000000852399949420;
	07: data <= 64'd0000001092647337676;
	08: data <= 64'd0000000852129179340;
	09: data <= 64'd0000000852129179340;
	10: data <= 64'd0000000852129179340;
	11: data <= 64'd0000000854276651894;
	12: data <= 64'd0000000000000000000;
	13: data <= 64'd0000000000000000000;
	14: data <= 64'd0000000000000000000;
	15: data <= 64'd0000000000000000000;
	//Alastal   
	16: data <= 64'd0000000000000000000;
	17: data <= 64'd0000000000000000000;
	18: data <= 64'd0075998244785848320;
	19: data <= 64'd0253890432214335488;
	20: data <= 64'd0488077612837601280;
	21: data <= 64'd0893534599569833984;
	22: data <= 64'd0893416474250674176;
	23: data <= 64'd1145740322541764608;
	24: data <= 64'd0893626360762826752;
	25: data <= 64'd0893625982805704704;
	26: data <= 64'd0893627580936192000;
	27: data <= 64'd0896065660304211968;
	28: data <= 64'd0000000000000000000;
	29: data <= 64'd0000000000000000000;
	30: data <= 64'd0000000000000000000;
	31: data <= 64'd0000000000000000000;
	default: data <= 64'b0;
	endcase
	end
endmodule 