// Original_Sine.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module Original_Sine (
		input  wire [14:0] a,      //      a.a
		input  wire        areset, // areset.reset
		output wire [13:0] c,      //      c.c
		input  wire        clk,    //    clk.clk
		output wire [13:0] s       //      s.s
	);

	Original_Sine_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.a      (a),      //      a.a
		.c      (c),      //      c.c
		.s      (s)       //      s.s
	);

endmodule
