// NiosII_Controlled_Section.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module NiosII_Controlled_Section (
		input  wire [7:0]  channel1_analog_export,     //     channel1_analog.export
		input  wire [7:0]  channel2_analog_export,     //     channel2_analog.export
		input  wire [7:0]  channel3_analog_export,     //     channel3_analog.export
		input  wire [7:0]  channel4_analog_export,     //     channel4_analog.export
		input  wire [7:0]  channel5_analog_export,     //     channel5_analog.export
		input  wire [7:0]  channel6_analog_export,     //     channel6_analog.export
		input  wire        clk_clk,                    //                 clk.clk
		output wire [11:0] read_address_export,        //        read_address.export
		input  wire        read_new_sample_export,     //     read_new_sample.export
		input  wire        reset_reset_n,              //               reset.reset_n
		inout  wire [15:0] sram_DQ,                    //                sram.DQ
		output wire [19:0] sram_ADDR,                  //                    .ADDR
		output wire        sram_LB_N,                  //                    .LB_N
		output wire        sram_UB_N,                  //                    .UB_N
		output wire        sram_CE_N,                  //                    .CE_N
		output wire        sram_OE_N,                  //                    .OE_N
		output wire        sram_WE_N,                  //                    .WE_N
		output wire        vga_CLK,                    //                 vga.CLK
		output wire        vga_HS,                     //                    .HS
		output wire        vga_VS,                     //                    .VS
		output wire        vga_BLANK,                  //                    .BLANK
		output wire        vga_SYNC,                   //                    .SYNC
		output wire [7:0]  vga_R,                      //                    .R
		output wire [7:0]  vga_G,                      //                    .G
		output wire [7:0]  vga_B,                      //                    .B
		output wire [10:1] H_Counter,
		output wire [10:1] V_Counter,
		input  wire        writing_finish_flag_export  // writing_finish_flag.export
	);

	wire         alpha_blender_avalon_blended_source_valid;                               // Alpha_Blender:output_valid -> FIFO:stream_in_valid
	wire  [29:0] alpha_blender_avalon_blended_source_data;                                // Alpha_Blender:output_data -> FIFO:stream_in_data
	wire         alpha_blender_avalon_blended_source_ready;                               // FIFO:stream_in_ready -> Alpha_Blender:output_ready
	wire         alpha_blender_avalon_blended_source_startofpacket;                       // Alpha_Blender:output_startofpacket -> FIFO:stream_in_startofpacket
	wire         alpha_blender_avalon_blended_source_endofpacket;                         // Alpha_Blender:output_endofpacket -> FIFO:stream_in_endofpacket
	wire         character_buffer_avalon_char_source_valid;                               // Character_Buffer:stream_valid -> Alpha_Blender:foreground_valid
	wire  [39:0] character_buffer_avalon_char_source_data;                                // Character_Buffer:stream_data -> Alpha_Blender:foreground_data
	wire         character_buffer_avalon_char_source_ready;                               // Alpha_Blender:foreground_ready -> Character_Buffer:stream_ready
	wire         character_buffer_avalon_char_source_startofpacket;                       // Character_Buffer:stream_startofpacket -> Alpha_Blender:foreground_startofpacket
	wire         character_buffer_avalon_char_source_endofpacket;                         // Character_Buffer:stream_endofpacket -> Alpha_Blender:foreground_endofpacket
	wire         fifo_avalon_dc_buffer_source_valid;                                      // FIFO:stream_out_valid -> VGA_Controller:valid
	wire  [29:0] fifo_avalon_dc_buffer_source_data;                                       // FIFO:stream_out_data -> VGA_Controller:data
	wire         fifo_avalon_dc_buffer_source_ready;                                      // VGA_Controller:ready -> FIFO:stream_out_ready
	wire         fifo_avalon_dc_buffer_source_startofpacket;                              // FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	wire         fifo_avalon_dc_buffer_source_endofpacket;                                // FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	wire         pixel_buffer_avalon_pixel_source_valid;                                  // Pixel_Buffer:stream_valid -> RGB_Resampler:stream_in_valid
	wire  [23:0] pixel_buffer_avalon_pixel_source_data;                                   // Pixel_Buffer:stream_data -> RGB_Resampler:stream_in_data
	wire         pixel_buffer_avalon_pixel_source_ready;                                  // RGB_Resampler:stream_in_ready -> Pixel_Buffer:stream_ready
	wire         pixel_buffer_avalon_pixel_source_startofpacket;                          // Pixel_Buffer:stream_startofpacket -> RGB_Resampler:stream_in_startofpacket
	wire         pixel_buffer_avalon_pixel_source_endofpacket;                            // Pixel_Buffer:stream_endofpacket -> RGB_Resampler:stream_in_endofpacket
	wire         rgb_resampler_avalon_rgb_source_valid;                                   // RGB_Resampler:stream_out_valid -> Alpha_Blender:background_valid
	wire  [29:0] rgb_resampler_avalon_rgb_source_data;                                    // RGB_Resampler:stream_out_data -> Alpha_Blender:background_data
	wire         rgb_resampler_avalon_rgb_source_ready;                                   // Alpha_Blender:background_ready -> RGB_Resampler:stream_out_ready
	wire         rgb_resampler_avalon_rgb_source_startofpacket;                           // RGB_Resampler:stream_out_startofpacket -> Alpha_Blender:background_startofpacket
	wire         rgb_resampler_avalon_rgb_source_endofpacket;                             // RGB_Resampler:stream_out_endofpacket -> Alpha_Blender:background_endofpacket
	wire         vga_pll_vga_clk_clk;                                                     // VGA_PLL:vga_clk_clk -> [FIFO:clk_stream_out, VGA_Controller:clk, rst_controller_001:clk]
	wire         pixel_buffer_avalon_pixel_dma_master_waitrequest;                        // mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_waitrequest -> Pixel_Buffer:master_waitrequest
	wire  [31:0] pixel_buffer_avalon_pixel_dma_master_readdata;                           // mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_readdata -> Pixel_Buffer:master_readdata
	wire  [31:0] pixel_buffer_avalon_pixel_dma_master_address;                            // Pixel_Buffer:master_address -> mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_address
	wire         pixel_buffer_avalon_pixel_dma_master_read;                               // Pixel_Buffer:master_read -> mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_read
	wire         pixel_buffer_avalon_pixel_dma_master_readdatavalid;                      // mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_readdatavalid -> Pixel_Buffer:master_readdatavalid
	wire         pixel_buffer_avalon_pixel_dma_master_lock;                               // Pixel_Buffer:master_arbiterlock -> mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_lock
	wire  [31:0] niosii_data_master_readdata;                                             // mm_interconnect_0:NiosII_data_master_readdata -> NiosII:d_readdata
	wire         niosii_data_master_waitrequest;                                          // mm_interconnect_0:NiosII_data_master_waitrequest -> NiosII:d_waitrequest
	wire         niosii_data_master_debugaccess;                                          // NiosII:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NiosII_data_master_debugaccess
	wire  [21:0] niosii_data_master_address;                                              // NiosII:d_address -> mm_interconnect_0:NiosII_data_master_address
	wire   [3:0] niosii_data_master_byteenable;                                           // NiosII:d_byteenable -> mm_interconnect_0:NiosII_data_master_byteenable
	wire         niosii_data_master_read;                                                 // NiosII:d_read -> mm_interconnect_0:NiosII_data_master_read
	wire         niosii_data_master_readdatavalid;                                        // mm_interconnect_0:NiosII_data_master_readdatavalid -> NiosII:d_readdatavalid
	wire         niosii_data_master_write;                                                // NiosII:d_write -> mm_interconnect_0:NiosII_data_master_write
	wire  [31:0] niosii_data_master_writedata;                                            // NiosII:d_writedata -> mm_interconnect_0:NiosII_data_master_writedata
	wire  [31:0] niosii_instruction_master_readdata;                                      // mm_interconnect_0:NiosII_instruction_master_readdata -> NiosII:i_readdata
	wire         niosii_instruction_master_waitrequest;                                   // mm_interconnect_0:NiosII_instruction_master_waitrequest -> NiosII:i_waitrequest
	wire  [21:0] niosii_instruction_master_address;                                       // NiosII:i_address -> mm_interconnect_0:NiosII_instruction_master_address
	wire         niosii_instruction_master_read;                                          // NiosII:i_read -> mm_interconnect_0:NiosII_instruction_master_read
	wire         niosii_instruction_master_readdatavalid;                                 // mm_interconnect_0:NiosII_instruction_master_readdatavalid -> NiosII:i_readdatavalid
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_readdata;                       // SRAM:readdata -> mm_interconnect_0:SRAM_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_avalon_sram_slave_address;                        // mm_interconnect_0:SRAM_avalon_sram_slave_address -> SRAM:address
	wire         mm_interconnect_0_sram_avalon_sram_slave_read;                           // mm_interconnect_0:SRAM_avalon_sram_slave_read -> SRAM:read
	wire   [1:0] mm_interconnect_0_sram_avalon_sram_slave_byteenable;                     // mm_interconnect_0:SRAM_avalon_sram_slave_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_avalon_sram_slave_readdatavalid;                  // SRAM:readdatavalid -> mm_interconnect_0:SRAM_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_avalon_sram_slave_write;                          // mm_interconnect_0:SRAM_avalon_sram_slave_write -> SRAM:write
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_writedata;                      // mm_interconnect_0:SRAM_avalon_sram_slave_writedata -> SRAM:writedata
	wire         mm_interconnect_0_character_buffer_avalon_char_buffer_slave_chipselect;  // mm_interconnect_0:Character_Buffer_avalon_char_buffer_slave_chipselect -> Character_Buffer:buf_chipselect
	wire   [7:0] mm_interconnect_0_character_buffer_avalon_char_buffer_slave_readdata;    // Character_Buffer:buf_readdata -> mm_interconnect_0:Character_Buffer_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_character_buffer_avalon_char_buffer_slave_waitrequest; // Character_Buffer:buf_waitrequest -> mm_interconnect_0:Character_Buffer_avalon_char_buffer_slave_waitrequest
	wire  [12:0] mm_interconnect_0_character_buffer_avalon_char_buffer_slave_address;     // mm_interconnect_0:Character_Buffer_avalon_char_buffer_slave_address -> Character_Buffer:buf_address
	wire         mm_interconnect_0_character_buffer_avalon_char_buffer_slave_read;        // mm_interconnect_0:Character_Buffer_avalon_char_buffer_slave_read -> Character_Buffer:buf_read
	wire   [0:0] mm_interconnect_0_character_buffer_avalon_char_buffer_slave_byteenable;  // mm_interconnect_0:Character_Buffer_avalon_char_buffer_slave_byteenable -> Character_Buffer:buf_byteenable
	wire         mm_interconnect_0_character_buffer_avalon_char_buffer_slave_write;       // mm_interconnect_0:Character_Buffer_avalon_char_buffer_slave_write -> Character_Buffer:buf_write
	wire   [7:0] mm_interconnect_0_character_buffer_avalon_char_buffer_slave_writedata;   // mm_interconnect_0:Character_Buffer_avalon_char_buffer_slave_writedata -> Character_Buffer:buf_writedata
	wire         mm_interconnect_0_character_buffer_avalon_char_control_slave_chipselect; // mm_interconnect_0:Character_Buffer_avalon_char_control_slave_chipselect -> Character_Buffer:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_character_buffer_avalon_char_control_slave_readdata;   // Character_Buffer:ctrl_readdata -> mm_interconnect_0:Character_Buffer_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_character_buffer_avalon_char_control_slave_address;    // mm_interconnect_0:Character_Buffer_avalon_char_control_slave_address -> Character_Buffer:ctrl_address
	wire         mm_interconnect_0_character_buffer_avalon_char_control_slave_read;       // mm_interconnect_0:Character_Buffer_avalon_char_control_slave_read -> Character_Buffer:ctrl_read
	wire   [3:0] mm_interconnect_0_character_buffer_avalon_char_control_slave_byteenable; // mm_interconnect_0:Character_Buffer_avalon_char_control_slave_byteenable -> Character_Buffer:ctrl_byteenable
	wire         mm_interconnect_0_character_buffer_avalon_char_control_slave_write;      // mm_interconnect_0:Character_Buffer_avalon_char_control_slave_write -> Character_Buffer:ctrl_write
	wire  [31:0] mm_interconnect_0_character_buffer_avalon_char_control_slave_writedata;  // mm_interconnect_0:Character_Buffer_avalon_char_control_slave_writedata -> Character_Buffer:ctrl_writedata
	wire  [31:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_readdata;            // Pixel_Buffer:slave_readdata -> mm_interconnect_0:Pixel_Buffer_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_address;             // mm_interconnect_0:Pixel_Buffer_avalon_control_slave_address -> Pixel_Buffer:slave_address
	wire         mm_interconnect_0_pixel_buffer_avalon_control_slave_read;                // mm_interconnect_0:Pixel_Buffer_avalon_control_slave_read -> Pixel_Buffer:slave_read
	wire   [3:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_byteenable;          // mm_interconnect_0:Pixel_Buffer_avalon_control_slave_byteenable -> Pixel_Buffer:slave_byteenable
	wire         mm_interconnect_0_pixel_buffer_avalon_control_slave_write;               // mm_interconnect_0:Pixel_Buffer_avalon_control_slave_write -> Pixel_Buffer:slave_write
	wire  [31:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_writedata;           // mm_interconnect_0:Pixel_Buffer_avalon_control_slave_writedata -> Pixel_Buffer:slave_writedata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                     // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                       // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                    // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                        // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                           // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                          // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                      // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire  [31:0] mm_interconnect_0_system_id_control_slave_readdata;                      // System_ID:readdata -> mm_interconnect_0:System_ID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_system_id_control_slave_address;                       // mm_interconnect_0:System_ID_control_slave_address -> System_ID:address
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_readdata;                       // NiosII:debug_mem_slave_readdata -> mm_interconnect_0:NiosII_debug_mem_slave_readdata
	wire         mm_interconnect_0_niosii_debug_mem_slave_waitrequest;                    // NiosII:debug_mem_slave_waitrequest -> mm_interconnect_0:NiosII_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_niosii_debug_mem_slave_debugaccess;                    // mm_interconnect_0:NiosII_debug_mem_slave_debugaccess -> NiosII:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_niosii_debug_mem_slave_address;                        // mm_interconnect_0:NiosII_debug_mem_slave_address -> NiosII:debug_mem_slave_address
	wire         mm_interconnect_0_niosii_debug_mem_slave_read;                           // mm_interconnect_0:NiosII_debug_mem_slave_read -> NiosII:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_niosii_debug_mem_slave_byteenable;                     // mm_interconnect_0:NiosII_debug_mem_slave_byteenable -> NiosII:debug_mem_slave_byteenable
	wire         mm_interconnect_0_niosii_debug_mem_slave_write;                          // mm_interconnect_0:NiosII_debug_mem_slave_write -> NiosII:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_writedata;                      // mm_interconnect_0:NiosII_debug_mem_slave_writedata -> NiosII:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                           // mm_interconnect_0:OnChip_Memory_s1_chipselect -> OnChip_Memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                             // OnChip_Memory:readdata -> mm_interconnect_0:OnChip_Memory_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory_s1_address;                              // mm_interconnect_0:OnChip_Memory_s1_address -> OnChip_Memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                           // mm_interconnect_0:OnChip_Memory_s1_byteenable -> OnChip_Memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                                // mm_interconnect_0:OnChip_Memory_s1_write -> OnChip_Memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                            // mm_interconnect_0:OnChip_Memory_s1_writedata -> OnChip_Memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                                // mm_interconnect_0:OnChip_Memory_s1_clken -> OnChip_Memory:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                                   // mm_interconnect_0:Timer_s1_chipselect -> Timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                     // Timer:readdata -> mm_interconnect_0:Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                      // mm_interconnect_0:Timer_s1_address -> Timer:address
	wire         mm_interconnect_0_timer_s1_write;                                        // mm_interconnect_0:Timer_s1_write -> Timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                                    // mm_interconnect_0:Timer_s1_writedata -> Timer:writedata
	wire  [31:0] mm_interconnect_0_channel1_analog_s1_readdata;                           // Channel1_Analog:readdata -> mm_interconnect_0:Channel1_Analog_s1_readdata
	wire   [1:0] mm_interconnect_0_channel1_analog_s1_address;                            // mm_interconnect_0:Channel1_Analog_s1_address -> Channel1_Analog:address
	wire  [31:0] mm_interconnect_0_channel2_analog_s1_readdata;                           // Channel2_Analog:readdata -> mm_interconnect_0:Channel2_Analog_s1_readdata
	wire   [1:0] mm_interconnect_0_channel2_analog_s1_address;                            // mm_interconnect_0:Channel2_Analog_s1_address -> Channel2_Analog:address
	wire  [31:0] mm_interconnect_0_channel3_analog_s1_readdata;                           // Channel3_Analog:readdata -> mm_interconnect_0:Channel3_Analog_s1_readdata
	wire   [1:0] mm_interconnect_0_channel3_analog_s1_address;                            // mm_interconnect_0:Channel3_Analog_s1_address -> Channel3_Analog:address
	wire  [31:0] mm_interconnect_0_channel4_analog_s1_readdata;                           // Channel4_Analog:readdata -> mm_interconnect_0:Channel4_Analog_s1_readdata
	wire   [1:0] mm_interconnect_0_channel4_analog_s1_address;                            // mm_interconnect_0:Channel4_Analog_s1_address -> Channel4_Analog:address
	wire  [31:0] mm_interconnect_0_channel5_analog_s1_readdata;                           // Channel5_Analog:readdata -> mm_interconnect_0:Channel5_Analog_s1_readdata
	wire   [1:0] mm_interconnect_0_channel5_analog_s1_address;                            // mm_interconnect_0:Channel5_Analog_s1_address -> Channel5_Analog:address
	wire  [31:0] mm_interconnect_0_channel6_analog_s1_readdata;                           // Channel6_Analog:readdata -> mm_interconnect_0:Channel6_Analog_s1_readdata
	wire   [1:0] mm_interconnect_0_channel6_analog_s1_address;                            // mm_interconnect_0:Channel6_Analog_s1_address -> Channel6_Analog:address
	wire  [31:0] mm_interconnect_0_writing_finish_flag_s1_readdata;                       // Writing_Finish_Flag:readdata -> mm_interconnect_0:Writing_Finish_Flag_s1_readdata
	wire   [1:0] mm_interconnect_0_writing_finish_flag_s1_address;                        // mm_interconnect_0:Writing_Finish_Flag_s1_address -> Writing_Finish_Flag:address
	wire  [31:0] mm_interconnect_0_read_new_sample_s1_readdata;                           // Read_New_Sample:readdata -> mm_interconnect_0:Read_New_Sample_s1_readdata
	wire   [1:0] mm_interconnect_0_read_new_sample_s1_address;                            // mm_interconnect_0:Read_New_Sample_s1_address -> Read_New_Sample:address
	wire         mm_interconnect_0_read_address_s1_chipselect;                            // mm_interconnect_0:Read_Address_s1_chipselect -> Read_Address:chipselect
	wire  [31:0] mm_interconnect_0_read_address_s1_readdata;                              // Read_Address:readdata -> mm_interconnect_0:Read_Address_s1_readdata
	wire   [1:0] mm_interconnect_0_read_address_s1_address;                               // mm_interconnect_0:Read_Address_s1_address -> Read_Address:address
	wire         mm_interconnect_0_read_address_s1_write;                                 // mm_interconnect_0:Read_Address_s1_write -> Read_Address:write_n
	wire  [31:0] mm_interconnect_0_read_address_s1_writedata;                             // mm_interconnect_0:Read_Address_s1_writedata -> Read_Address:writedata
	wire         irq_mapper_receiver0_irq;                                                // JTAG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                // Timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] niosii_irq_irq;                                                          // irq_mapper:sender_irq -> NiosII:irq
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [Alpha_Blender:reset, Channel1_Analog:reset_n, Channel2_Analog:reset_n, Channel3_Analog:reset_n, Channel4_Analog:reset_n, Channel5_Analog:reset_n, Channel6_Analog:reset_n, Character_Buffer:reset, FIFO:reset_stream_in, JTAG:rst_n, NiosII:reset_n, OnChip_Memory:reset, Pixel_Buffer:reset, RGB_Resampler:reset, Read_Address:reset_n, Read_New_Sample:reset_n, SRAM:reset, System_ID:reset_n, Timer:reset_n, VGA_PLL:ref_reset_reset, Writing_Finish_Flag:reset_n, irq_mapper:reset, mm_interconnect_0:Pixel_Buffer_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [NiosII:reset_req, OnChip_Memory:reset_req, rst_translator:reset_req_in]
	wire         niosii_debug_reset_request_reset;                                        // NiosII:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         vga_pll_reset_source_reset;                                              // VGA_PLL:reset_source_reset -> [rst_controller:reset_in2, rst_controller_001:reset_in2]
	wire         rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> [FIFO:reset_stream_out, VGA_Controller:reset]

	NiosII_Controlled_Section_Alpha_Blender alpha_blender (
		.clk                      (clk_clk),                                           //                    clk.clk
		.reset                    (rst_controller_reset_out_reset),                    //                  reset.reset
		.foreground_data          (character_buffer_avalon_char_source_data),          // avalon_foreground_sink.data
		.foreground_startofpacket (character_buffer_avalon_char_source_startofpacket), //                       .startofpacket
		.foreground_endofpacket   (character_buffer_avalon_char_source_endofpacket),   //                       .endofpacket
		.foreground_valid         (character_buffer_avalon_char_source_valid),         //                       .valid
		.foreground_ready         (character_buffer_avalon_char_source_ready),         //                       .ready
		.background_data          (rgb_resampler_avalon_rgb_source_data),              // avalon_background_sink.data
		.background_startofpacket (rgb_resampler_avalon_rgb_source_startofpacket),     //                       .startofpacket
		.background_endofpacket   (rgb_resampler_avalon_rgb_source_endofpacket),       //                       .endofpacket
		.background_valid         (rgb_resampler_avalon_rgb_source_valid),             //                       .valid
		.background_ready         (rgb_resampler_avalon_rgb_source_ready),             //                       .ready
		.output_ready             (alpha_blender_avalon_blended_source_ready),         //  avalon_blended_source.ready
		.output_data              (alpha_blender_avalon_blended_source_data),          //                       .data
		.output_startofpacket     (alpha_blender_avalon_blended_source_startofpacket), //                       .startofpacket
		.output_endofpacket       (alpha_blender_avalon_blended_source_endofpacket),   //                       .endofpacket
		.output_valid             (alpha_blender_avalon_blended_source_valid)          //                       .valid
	);

	NiosII_Controlled_Section_Channel1_Analog channel1_analog (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_channel1_analog_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_channel1_analog_s1_readdata), //                    .readdata
		.in_port  (channel1_analog_export)                         // external_connection.export
	);

	NiosII_Controlled_Section_Channel1_Analog channel2_analog (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_channel2_analog_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_channel2_analog_s1_readdata), //                    .readdata
		.in_port  (channel2_analog_export)                         // external_connection.export
	);

	NiosII_Controlled_Section_Channel1_Analog channel3_analog (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_channel3_analog_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_channel3_analog_s1_readdata), //                    .readdata
		.in_port  (channel3_analog_export)                         // external_connection.export
	);

	NiosII_Controlled_Section_Channel1_Analog channel4_analog (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_channel4_analog_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_channel4_analog_s1_readdata), //                    .readdata
		.in_port  (channel4_analog_export)                         // external_connection.export
	);

	NiosII_Controlled_Section_Channel1_Analog channel5_analog (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_channel5_analog_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_channel5_analog_s1_readdata), //                    .readdata
		.in_port  (channel5_analog_export)                         // external_connection.export
	);

	NiosII_Controlled_Section_Channel1_Analog channel6_analog (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_channel6_analog_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_channel6_analog_s1_readdata), //                    .readdata
		.in_port  (channel6_analog_export)                         // external_connection.export
	);

	NiosII_Controlled_Section_Character_Buffer character_buffer (
		.clk                  (clk_clk),                                                                 //                       clk.clk
		.reset                (rst_controller_reset_out_reset),                                          //                     reset.reset
		.ctrl_address         (mm_interconnect_0_character_buffer_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_character_buffer_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_character_buffer_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_character_buffer_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_character_buffer_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_character_buffer_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_character_buffer_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (character_buffer_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (character_buffer_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (character_buffer_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (character_buffer_avalon_char_source_valid),                               //                          .valid
		.stream_data          (character_buffer_avalon_char_source_data)                                 //                          .data
	);

	NiosII_Controlled_Section_FIFO fifo (
		.clk_stream_in            (clk_clk),                                           //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                    //         reset_stream_in.reset
		.clk_stream_out           (vga_pll_vga_clk_clk),                               //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_001_reset_out_reset),                //        reset_stream_out.reset
		.stream_in_ready          (alpha_blender_avalon_blended_source_ready),         //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (alpha_blender_avalon_blended_source_startofpacket), //                        .startofpacket
		.stream_in_endofpacket    (alpha_blender_avalon_blended_source_endofpacket),   //                        .endofpacket
		.stream_in_valid          (alpha_blender_avalon_blended_source_valid),         //                        .valid
		.stream_in_data           (alpha_blender_avalon_blended_source_data),          //                        .data
		.stream_out_ready         (fifo_avalon_dc_buffer_source_ready),                // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (fifo_avalon_dc_buffer_source_startofpacket),        //                        .startofpacket
		.stream_out_endofpacket   (fifo_avalon_dc_buffer_source_endofpacket),          //                        .endofpacket
		.stream_out_valid         (fifo_avalon_dc_buffer_source_valid),                //                        .valid
		.stream_out_data          (fifo_avalon_dc_buffer_source_data)                  //                        .data
	);

	NiosII_Controlled_Section_JTAG jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	NiosII_Controlled_Section_NiosII niosii (
		.clk                                 (clk_clk),                                              //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (niosii_data_master_address),                           //               data_master.address
		.d_byteenable                        (niosii_data_master_byteenable),                        //                          .byteenable
		.d_read                              (niosii_data_master_read),                              //                          .read
		.d_readdata                          (niosii_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (niosii_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (niosii_data_master_write),                             //                          .write
		.d_writedata                         (niosii_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (niosii_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (niosii_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (niosii_instruction_master_address),                    //        instruction_master.address
		.i_read                              (niosii_instruction_master_read),                       //                          .read
		.i_readdata                          (niosii_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (niosii_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (niosii_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (niosii_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (niosii_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_niosii_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_niosii_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_niosii_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_niosii_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_niosii_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_niosii_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_niosii_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_niosii_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	NiosII_Controlled_Section_OnChip_Memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	NiosII_Controlled_Section_Pixel_Buffer pixel_buffer (
		.clk                  (clk_clk),                                                        //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                                 //                   reset.reset
		.master_readdatavalid (pixel_buffer_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (pixel_buffer_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (pixel_buffer_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (pixel_buffer_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (pixel_buffer_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_pixel_buffer_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_pixel_buffer_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_pixel_buffer_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_pixel_buffer_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_pixel_buffer_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_pixel_buffer_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (pixel_buffer_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (pixel_buffer_avalon_pixel_source_data)                           //                        .data
	);

	NiosII_Controlled_Section_RGB_Resampler rgb_resampler (
		.clk                      (clk_clk),                                        //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                 //             reset.reset
		.stream_in_startofpacket  (pixel_buffer_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (pixel_buffer_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (pixel_buffer_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (pixel_buffer_avalon_pixel_source_data),          //                  .data
		.slave_read               (),                                               //  avalon_rgb_slave.read
		.slave_readdata           (),                                               //                  .readdata
		.stream_out_ready         (rgb_resampler_avalon_rgb_source_ready),          // avalon_rgb_source.ready
		.stream_out_startofpacket (rgb_resampler_avalon_rgb_source_startofpacket),  //                  .startofpacket
		.stream_out_endofpacket   (rgb_resampler_avalon_rgb_source_endofpacket),    //                  .endofpacket
		.stream_out_valid         (rgb_resampler_avalon_rgb_source_valid),          //                  .valid
		.stream_out_data          (rgb_resampler_avalon_rgb_source_data)            //                  .data
	);

	NiosII_Controlled_Section_Read_Address read_address (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_read_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_read_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_read_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_read_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_read_address_s1_readdata),   //                    .readdata
		.out_port   (read_address_export)                           // external_connection.export
	);

	NiosII_Controlled_Section_Read_New_Sample read_new_sample (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_read_new_sample_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_read_new_sample_s1_readdata), //                    .readdata
		.in_port  (read_new_sample_export)                         // external_connection.export
	);

	NiosII_Controlled_Section_SRAM sram (
		.clk           (clk_clk),                                                //                clk.clk
		.reset         (rst_controller_reset_out_reset),                         //              reset.reset
		.SRAM_DQ       (sram_DQ),                                                // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                              //                   .export
		.SRAM_LB_N     (sram_LB_N),                                              //                   .export
		.SRAM_UB_N     (sram_UB_N),                                              //                   .export
		.SRAM_CE_N     (sram_CE_N),                                              //                   .export
		.SRAM_OE_N     (sram_OE_N),                                              //                   .export
		.SRAM_WE_N     (sram_WE_N),                                              //                   .export
		.address       (mm_interconnect_0_sram_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	NiosII_Controlled_Section_System_ID system_id (
		.clock    (clk_clk),                                            //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                    //         reset.reset_n
		.readdata (mm_interconnect_0_system_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_system_id_control_slave_address)   //              .address
	);

	NiosII_Controlled_Section_Timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	NiosII_Controlled_Section_VGA_Controller vga_controller (
		.clk           (vga_pll_vga_clk_clk),                        //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),         //              reset.reset
		.data          (fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_CLK),                                    // external_interface.export
		.VGA_HS        (vga_HS),                                     //                   .export
		.VGA_VS        (vga_VS),                                     //                   .export
		.VGA_BLANK     (vga_BLANK),                                  //                   .export
		.VGA_SYNC      (vga_SYNC),                                   //                   .export
		.H_Counter		(H_Counter),
		.V_Counter		(V_Counter),
		.VGA_R         (vga_R),                                      //                   .export
		.VGA_G         (vga_G),                                      //                   .export
		.VGA_B         (vga_B)                                       //                   .export
	);

	NiosII_Controlled_Section_VGA_PLL vga_pll (
		.ref_clk_clk        (clk_clk),                        //      ref_clk.clk
		.ref_reset_reset    (rst_controller_reset_out_reset), //    ref_reset.reset
		.vga_clk_clk        (vga_pll_vga_clk_clk),            //      vga_clk.clk
		.reset_source_reset (vga_pll_reset_source_reset)      // reset_source.reset
	);

	NiosII_Controlled_Section_Read_New_Sample writing_finish_flag (
		.clk      (clk_clk),                                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (mm_interconnect_0_writing_finish_flag_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_writing_finish_flag_s1_readdata), //                    .readdata
		.in_port  (writing_finish_flag_export)                         // external_connection.export
	);

	NiosII_Controlled_Section_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                         (clk_clk),                                                                 //                                  clk_0_clk.clk
		.Pixel_Buffer_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                                          //   Pixel_Buffer_reset_reset_bridge_in_reset.reset
		.NiosII_data_master_address                            (niosii_data_master_address),                                              //                         NiosII_data_master.address
		.NiosII_data_master_waitrequest                        (niosii_data_master_waitrequest),                                          //                                           .waitrequest
		.NiosII_data_master_byteenable                         (niosii_data_master_byteenable),                                           //                                           .byteenable
		.NiosII_data_master_read                               (niosii_data_master_read),                                                 //                                           .read
		.NiosII_data_master_readdata                           (niosii_data_master_readdata),                                             //                                           .readdata
		.NiosII_data_master_readdatavalid                      (niosii_data_master_readdatavalid),                                        //                                           .readdatavalid
		.NiosII_data_master_write                              (niosii_data_master_write),                                                //                                           .write
		.NiosII_data_master_writedata                          (niosii_data_master_writedata),                                            //                                           .writedata
		.NiosII_data_master_debugaccess                        (niosii_data_master_debugaccess),                                          //                                           .debugaccess
		.NiosII_instruction_master_address                     (niosii_instruction_master_address),                                       //                  NiosII_instruction_master.address
		.NiosII_instruction_master_waitrequest                 (niosii_instruction_master_waitrequest),                                   //                                           .waitrequest
		.NiosII_instruction_master_read                        (niosii_instruction_master_read),                                          //                                           .read
		.NiosII_instruction_master_readdata                    (niosii_instruction_master_readdata),                                      //                                           .readdata
		.NiosII_instruction_master_readdatavalid               (niosii_instruction_master_readdatavalid),                                 //                                           .readdatavalid
		.Pixel_Buffer_avalon_pixel_dma_master_address          (pixel_buffer_avalon_pixel_dma_master_address),                            //       Pixel_Buffer_avalon_pixel_dma_master.address
		.Pixel_Buffer_avalon_pixel_dma_master_waitrequest      (pixel_buffer_avalon_pixel_dma_master_waitrequest),                        //                                           .waitrequest
		.Pixel_Buffer_avalon_pixel_dma_master_read             (pixel_buffer_avalon_pixel_dma_master_read),                               //                                           .read
		.Pixel_Buffer_avalon_pixel_dma_master_readdata         (pixel_buffer_avalon_pixel_dma_master_readdata),                           //                                           .readdata
		.Pixel_Buffer_avalon_pixel_dma_master_readdatavalid    (pixel_buffer_avalon_pixel_dma_master_readdatavalid),                      //                                           .readdatavalid
		.Pixel_Buffer_avalon_pixel_dma_master_lock             (pixel_buffer_avalon_pixel_dma_master_lock),                               //                                           .lock
		.Channel1_Analog_s1_address                            (mm_interconnect_0_channel1_analog_s1_address),                            //                         Channel1_Analog_s1.address
		.Channel1_Analog_s1_readdata                           (mm_interconnect_0_channel1_analog_s1_readdata),                           //                                           .readdata
		.Channel2_Analog_s1_address                            (mm_interconnect_0_channel2_analog_s1_address),                            //                         Channel2_Analog_s1.address
		.Channel2_Analog_s1_readdata                           (mm_interconnect_0_channel2_analog_s1_readdata),                           //                                           .readdata
		.Channel3_Analog_s1_address                            (mm_interconnect_0_channel3_analog_s1_address),                            //                         Channel3_Analog_s1.address
		.Channel3_Analog_s1_readdata                           (mm_interconnect_0_channel3_analog_s1_readdata),                           //                                           .readdata
		.Channel4_Analog_s1_address                            (mm_interconnect_0_channel4_analog_s1_address),                            //                         Channel4_Analog_s1.address
		.Channel4_Analog_s1_readdata                           (mm_interconnect_0_channel4_analog_s1_readdata),                           //                                           .readdata
		.Channel5_Analog_s1_address                            (mm_interconnect_0_channel5_analog_s1_address),                            //                         Channel5_Analog_s1.address
		.Channel5_Analog_s1_readdata                           (mm_interconnect_0_channel5_analog_s1_readdata),                           //                                           .readdata
		.Channel6_Analog_s1_address                            (mm_interconnect_0_channel6_analog_s1_address),                            //                         Channel6_Analog_s1.address
		.Channel6_Analog_s1_readdata                           (mm_interconnect_0_channel6_analog_s1_readdata),                           //                                           .readdata
		.Character_Buffer_avalon_char_buffer_slave_address     (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_address),     //  Character_Buffer_avalon_char_buffer_slave.address
		.Character_Buffer_avalon_char_buffer_slave_write       (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_write),       //                                           .write
		.Character_Buffer_avalon_char_buffer_slave_read        (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_read),        //                                           .read
		.Character_Buffer_avalon_char_buffer_slave_readdata    (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_readdata),    //                                           .readdata
		.Character_Buffer_avalon_char_buffer_slave_writedata   (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_writedata),   //                                           .writedata
		.Character_Buffer_avalon_char_buffer_slave_byteenable  (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_byteenable),  //                                           .byteenable
		.Character_Buffer_avalon_char_buffer_slave_waitrequest (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_waitrequest), //                                           .waitrequest
		.Character_Buffer_avalon_char_buffer_slave_chipselect  (mm_interconnect_0_character_buffer_avalon_char_buffer_slave_chipselect),  //                                           .chipselect
		.Character_Buffer_avalon_char_control_slave_address    (mm_interconnect_0_character_buffer_avalon_char_control_slave_address),    // Character_Buffer_avalon_char_control_slave.address
		.Character_Buffer_avalon_char_control_slave_write      (mm_interconnect_0_character_buffer_avalon_char_control_slave_write),      //                                           .write
		.Character_Buffer_avalon_char_control_slave_read       (mm_interconnect_0_character_buffer_avalon_char_control_slave_read),       //                                           .read
		.Character_Buffer_avalon_char_control_slave_readdata   (mm_interconnect_0_character_buffer_avalon_char_control_slave_readdata),   //                                           .readdata
		.Character_Buffer_avalon_char_control_slave_writedata  (mm_interconnect_0_character_buffer_avalon_char_control_slave_writedata),  //                                           .writedata
		.Character_Buffer_avalon_char_control_slave_byteenable (mm_interconnect_0_character_buffer_avalon_char_control_slave_byteenable), //                                           .byteenable
		.Character_Buffer_avalon_char_control_slave_chipselect (mm_interconnect_0_character_buffer_avalon_char_control_slave_chipselect), //                                           .chipselect
		.JTAG_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_avalon_jtag_slave_address),                        //                     JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_avalon_jtag_slave_write),                          //                                           .write
		.JTAG_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_avalon_jtag_slave_read),                           //                                           .read
		.JTAG_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                       //                                           .readdata
		.JTAG_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),                      //                                           .writedata
		.JTAG_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),                    //                                           .waitrequest
		.JTAG_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),                     //                                           .chipselect
		.NiosII_debug_mem_slave_address                        (mm_interconnect_0_niosii_debug_mem_slave_address),                        //                     NiosII_debug_mem_slave.address
		.NiosII_debug_mem_slave_write                          (mm_interconnect_0_niosii_debug_mem_slave_write),                          //                                           .write
		.NiosII_debug_mem_slave_read                           (mm_interconnect_0_niosii_debug_mem_slave_read),                           //                                           .read
		.NiosII_debug_mem_slave_readdata                       (mm_interconnect_0_niosii_debug_mem_slave_readdata),                       //                                           .readdata
		.NiosII_debug_mem_slave_writedata                      (mm_interconnect_0_niosii_debug_mem_slave_writedata),                      //                                           .writedata
		.NiosII_debug_mem_slave_byteenable                     (mm_interconnect_0_niosii_debug_mem_slave_byteenable),                     //                                           .byteenable
		.NiosII_debug_mem_slave_waitrequest                    (mm_interconnect_0_niosii_debug_mem_slave_waitrequest),                    //                                           .waitrequest
		.NiosII_debug_mem_slave_debugaccess                    (mm_interconnect_0_niosii_debug_mem_slave_debugaccess),                    //                                           .debugaccess
		.OnChip_Memory_s1_address                              (mm_interconnect_0_onchip_memory_s1_address),                              //                           OnChip_Memory_s1.address
		.OnChip_Memory_s1_write                                (mm_interconnect_0_onchip_memory_s1_write),                                //                                           .write
		.OnChip_Memory_s1_readdata                             (mm_interconnect_0_onchip_memory_s1_readdata),                             //                                           .readdata
		.OnChip_Memory_s1_writedata                            (mm_interconnect_0_onchip_memory_s1_writedata),                            //                                           .writedata
		.OnChip_Memory_s1_byteenable                           (mm_interconnect_0_onchip_memory_s1_byteenable),                           //                                           .byteenable
		.OnChip_Memory_s1_chipselect                           (mm_interconnect_0_onchip_memory_s1_chipselect),                           //                                           .chipselect
		.OnChip_Memory_s1_clken                                (mm_interconnect_0_onchip_memory_s1_clken),                                //                                           .clken
		.Pixel_Buffer_avalon_control_slave_address             (mm_interconnect_0_pixel_buffer_avalon_control_slave_address),             //          Pixel_Buffer_avalon_control_slave.address
		.Pixel_Buffer_avalon_control_slave_write               (mm_interconnect_0_pixel_buffer_avalon_control_slave_write),               //                                           .write
		.Pixel_Buffer_avalon_control_slave_read                (mm_interconnect_0_pixel_buffer_avalon_control_slave_read),                //                                           .read
		.Pixel_Buffer_avalon_control_slave_readdata            (mm_interconnect_0_pixel_buffer_avalon_control_slave_readdata),            //                                           .readdata
		.Pixel_Buffer_avalon_control_slave_writedata           (mm_interconnect_0_pixel_buffer_avalon_control_slave_writedata),           //                                           .writedata
		.Pixel_Buffer_avalon_control_slave_byteenable          (mm_interconnect_0_pixel_buffer_avalon_control_slave_byteenable),          //                                           .byteenable
		.Read_Address_s1_address                               (mm_interconnect_0_read_address_s1_address),                               //                            Read_Address_s1.address
		.Read_Address_s1_write                                 (mm_interconnect_0_read_address_s1_write),                                 //                                           .write
		.Read_Address_s1_readdata                              (mm_interconnect_0_read_address_s1_readdata),                              //                                           .readdata
		.Read_Address_s1_writedata                             (mm_interconnect_0_read_address_s1_writedata),                             //                                           .writedata
		.Read_Address_s1_chipselect                            (mm_interconnect_0_read_address_s1_chipselect),                            //                                           .chipselect
		.Read_New_Sample_s1_address                            (mm_interconnect_0_read_new_sample_s1_address),                            //                         Read_New_Sample_s1.address
		.Read_New_Sample_s1_readdata                           (mm_interconnect_0_read_new_sample_s1_readdata),                           //                                           .readdata
		.SRAM_avalon_sram_slave_address                        (mm_interconnect_0_sram_avalon_sram_slave_address),                        //                     SRAM_avalon_sram_slave.address
		.SRAM_avalon_sram_slave_write                          (mm_interconnect_0_sram_avalon_sram_slave_write),                          //                                           .write
		.SRAM_avalon_sram_slave_read                           (mm_interconnect_0_sram_avalon_sram_slave_read),                           //                                           .read
		.SRAM_avalon_sram_slave_readdata                       (mm_interconnect_0_sram_avalon_sram_slave_readdata),                       //                                           .readdata
		.SRAM_avalon_sram_slave_writedata                      (mm_interconnect_0_sram_avalon_sram_slave_writedata),                      //                                           .writedata
		.SRAM_avalon_sram_slave_byteenable                     (mm_interconnect_0_sram_avalon_sram_slave_byteenable),                     //                                           .byteenable
		.SRAM_avalon_sram_slave_readdatavalid                  (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid),                  //                                           .readdatavalid
		.System_ID_control_slave_address                       (mm_interconnect_0_system_id_control_slave_address),                       //                    System_ID_control_slave.address
		.System_ID_control_slave_readdata                      (mm_interconnect_0_system_id_control_slave_readdata),                      //                                           .readdata
		.Timer_s1_address                                      (mm_interconnect_0_timer_s1_address),                                      //                                   Timer_s1.address
		.Timer_s1_write                                        (mm_interconnect_0_timer_s1_write),                                        //                                           .write
		.Timer_s1_readdata                                     (mm_interconnect_0_timer_s1_readdata),                                     //                                           .readdata
		.Timer_s1_writedata                                    (mm_interconnect_0_timer_s1_writedata),                                    //                                           .writedata
		.Timer_s1_chipselect                                   (mm_interconnect_0_timer_s1_chipselect),                                   //                                           .chipselect
		.Writing_Finish_Flag_s1_address                        (mm_interconnect_0_writing_finish_flag_s1_address),                        //                     Writing_Finish_Flag_s1.address
		.Writing_Finish_Flag_s1_readdata                       (mm_interconnect_0_writing_finish_flag_s1_readdata)                        //                                           .readdata
	);

	NiosII_Controlled_Section_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (niosii_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (niosii_debug_reset_request_reset),   // reset_in1.reset
		.reset_in2      (vga_pll_reset_source_reset),         // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (niosii_debug_reset_request_reset),   // reset_in1.reset
		.reset_in2      (vga_pll_reset_source_reset),         // reset_in2.reset
		.clk            (vga_pll_vga_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
