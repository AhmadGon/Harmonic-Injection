module HarmonicROM(
	input VGA_CLK,
	input [5:0] address,
	output reg [31:0] data
);
always @(posedge VGA_CLK)
	begin
	case(address)
	//M
	00: data <= 32'b00000000000000000000000000000000;
	01: data <= 32'b00000000000000000000000000000000;
	02: data <= 32'b11000011000000000000000000000000;
	03: data <= 32'b11100111000000000000000000000000;
	04: data <= 32'b11111111000000000000000000000000;
	05: data <= 32'b11111111000000000000000000000000;
	06: data <= 32'b11011011000000000000000000000000;
	07: data <= 32'b11000011000000000000000000000000;
	08: data <= 32'b11000011000000000000000000000000;
	09: data <= 32'b11000011000000000000000000000000;
	10: data <= 32'b11000011000000000000000000000000;
	11: data <= 32'b11000011000000000000000000000000;
	12: data <= 32'b00000000000000000000000000000000;
	13: data <= 32'b00000000000000000000000000000000;
	14: data <= 32'b00000000000000000000000000000000;
	15: data <= 32'b00000000000000000000000000000000;
	//3rd 
	16: data <= 32'b00000000000000000000000000000000;
	17: data <= 32'b00000000000000000000000000000000;
	18: data <= 32'b01111100000000000001110000000000;
	19: data <= 32'b11000110000000000000110000000000;
	20: data <= 32'b00000110000000000000110000000000;
	21: data <= 32'b00000110110111000011110000000000;
	22: data <= 32'b00111100011101100110110000000000;
	23: data <= 32'b00000110011001101100110000000000;
	24: data <= 32'b00000110011000001100110000000000;
	25: data <= 32'b00000110011000001100110000000000;
	26: data <= 32'b11000110011000001100110000000000;
	27: data <= 32'b01111100111100000111011000000000;
	28: data <= 32'b00000000000000000000000000000000;
	29: data <= 32'b00000000000000000000000000000000;
	30: data <= 32'b00000000000000000000000000000000;
	31: data <= 32'b00000000000000000000000000000000;
	//9th
	32: data <= 32'b00000000000000000000000000000000;
	33: data <= 32'b00000000000000000000000000000000;
	34: data <= 32'b01111100000100001110000000000000;
	35: data <= 32'b11000110001100000110000000000000;
	36: data <= 32'b11000110001100000110000000000000;
	37: data <= 32'b11000110111111000110110000000000;
	38: data <= 32'b01111110001100000111011000000000;
	39: data <= 32'b00000110001100000110011000000000;
	40: data <= 32'b00000110001100000110011000000000;
	41: data <= 32'b00000110001100000110011000000000;
	42: data <= 32'b00001100001101100110011000000000;
	43: data <= 32'b01111000000111001110011000000000;
	44: data <= 32'b00000000000000000000000000000000;
	45: data <= 32'b00000000000000000000000000000000;
	46: data <= 32'b00000000000000000000000000000000;
	47: data <= 32'b00000000000000000000000000000000;
	//15th
	48: data <= 32'b00000000000000000000000000000000;
	49: data <= 32'b00000000000000000000000000000000;
	50: data <= 32'b00011000111111100001000011100000;
	51: data <= 32'b00111000110000000011000001100000;
	52: data <= 32'b01111000110000000011000001100000;
	53: data <= 32'b00011000110000001111110001101100;
	54: data <= 32'b00011000111111000011000001110110;
	55: data <= 32'b00011000000001100011000001100110;
	56: data <= 32'b00011000000001100011000001100110;
	57: data <= 32'b00011000000001100011000001100110;
	58: data <= 32'b00011000110001100011011001100110;
	59: data <= 32'b01111110011111000001110011100110;
	60: data <= 32'b00000000000000000000000000000000;
	61: data <= 32'b00000000000000000000000000000000;
	62: data <= 32'b00000000000000000000000000000000;
	63: data <= 32'b00000000000000000000000000000000;
	default: data <= 64'b0;
	endcase
	end
endmodule 