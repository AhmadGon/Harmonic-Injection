module StringROM(
	input VGA_CLK,
	input [5:0] address,
	output reg [63:0] data
);

always @(posedge VGA_CLK)
	begin
	case(address)
	//Phase A
	00: data <= 64'b0000000111111111111111111111111111111111111111111111111100000000;
	01: data <= 64'b0000011111111111111111111111111111111111111111111111111111000000;
	02: data <= 64'b0000011000000000000000000000000000000000000000000000000011000000;
	03: data <= 64'b0000110011111100111000000000000000000000000000000001000001100000;
	04: data <= 64'b0000110001100110011000000000000000000000000000000011100001100000;
	05: data <= 64'b0001100001100110011000000000000000000000000000000110110000110000;
	06: data <= 64'b0001100001100110011011000111100001111100011111001100011000110000;
	07: data <= 64'b0001100001111100011101100000110011000110110001101100011000110000;
	08: data <= 64'b0001100001100000011001100111110001100000111111101111111000110000;
	09: data <= 64'b0001100001100000011001101100110000111000110000001100011000110000;
	10: data <= 64'b0001100001100000011001101100110000001100110000001100011000110000;
	11: data <= 64'b0000110001100000011001101100110011000110110001101100011001100000;
	12: data <= 64'b0000110011110000111001100111011001111100011111001100011001100000;
	13: data <= 64'b0000011000000000000000000000000000000000000000000000000011000000;
	14: data <= 64'b0000011111111111111111111111111111111111111111111111111111000000;
	15: data <= 64'b0000000111111111111111111111111111111111111111111111111100000000;
	//Phase B   
	16: data <= 64'b0000000111111111111111111111111111111111111111111111111100000000;
	17: data <= 64'b0000011111111111111111111111111111111111111111111111111111000000;
	18: data <= 64'b0000011000000000000000000000000000000000000000000000000011000000;
	19: data <= 64'b0000110011111100111000000000000000000000000000001111110001100000;
	20: data <= 64'b0000110001100110011000000000000000000000000000000110011001100000;
	21: data <= 64'b0001100001100110011000000000000000000000000000000110011000110000;
	22: data <= 64'b0001100001100110011011000111100001111100011111000110011000110000;
	23: data <= 64'b0001100001111100011101100000110011000110110001100111110000110000;
	24: data <= 64'b0001100001100000011001100111110001100000111111100110011000110000;
	25: data <= 64'b0001100001100000011001101100110000111000110000000110011000110000;
	26: data <= 64'b0001100001100000011001101100110000001100110000000110011000110000;
	27: data <= 64'b0000110001100000011001101100110011000110110001100110011001100000;
	28: data <= 64'b0000110011110000111001100111011001111100011111001111110001100000;
	29: data <= 64'b0000011000000000000000000000000000000000000000000000000011000000;
	30: data <= 64'b0000011111111111111111111111111111111111111111111111111111000000;
	31: data <= 64'b0000000111111111111111111111111111111111111111111111111100000000;
	//Phase C
	32: data <= 64'b0000000111111111111111111111111111111111111111111111111100000000;
	33: data <= 64'b0000011111111111111111111111111111111111111111111111111111000000;
	34: data <= 64'b0000011000000000000000000000000000000000000000000000000011000000;
	35: data <= 64'b0000110011111100111000000000000000000000000000000011110001100000;
	36: data <= 64'b0000110001100110011000000000000000000000000000000110011001100000;
	37: data <= 64'b0001100001100110011000000000000000000000000000001100001000110000;
	38: data <= 64'b0001100001100110011011000111100001111100011111001100000000110000;
	39: data <= 64'b0001100001111100011101100000110011000110110001101100000000110000;
	40: data <= 64'b0001100001100000011001100111110001100000111111101100000000110000;
	41: data <= 64'b0001100001100000011001101100110000111000110000001100000000110000;
	42: data <= 64'b0001100001100000011001101100110000001100110000001100001000110000;
	43: data <= 64'b0000110001100000011001101100110011000110110001100110011001100000;
	44: data <= 64'b0000110011110000111001100111011001111100011111000011110001100000;
	45: data <= 64'b0000011000000000000000000000000000000000000000000000000011000000;
	46: data <= 64'b0000011111111111111111111111111111111111111111111111111111000000;
	47: data <= 64'b0000000111111111111111111111111111111111111111111111111100000000;
	default: data <= 64'b0;
	endcase
	end
endmodule 