
module Original_Sine (
	clk,
	areset,
	a,
	c,
	s);	

	input		clk;
	input		areset;
	input	[14:0]	a;
	output	[13:0]	c;
	output	[13:0]	s;
endmodule
